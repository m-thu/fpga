-- UART RX (9600, N, 8, 1)

-- ghdl -a --std=08 baudrate_gen.vhd
-- ghdl -a --std=08 uart_rx.vhd

-- Oversampling factor: 16
--
-- ------|    |----|    |- ... |----|----
--       |    |    |    |      |
--       |    |    |    |      |
--       |____|    |____|      |
-- idle   start d0   d1    ...  stop idle
--       ^  ^    ^
--       |  |    |
--       |  |    --- sample = 15, reset to 0
--       |  -------- sample =  7, reset to 0
--       ----------- sample =  0
--
-- IDLE  |START| DATA          | STOP     (FSM states)

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity uart_rx is
	port (
		clk, rst : in std_logic;
		rx : in std_logic;
		-- Gets asserted for one clock cycle when data is valid
		done : out std_logic;
		data : out std_logic_vector (7 downto 0)
	);
end entity;

architecture behav of uart_rx is
	type state_type is (IDLE, START, RDATA, STOP);
	signal tick : std_logic;
	signal state, next_state : state_type;
	
	-- Current data bit
	signal n, next_n : unsigned (2 downto 0);
	-- Received data
	signal rx_data, next_rx_data : std_logic_vector (7 downto 0);
	-- Sampling counter
	signal sample_count, next_sample_count : unsigned (3 downto 0);
begin
	-- Baudrate: 9600
	baudrate_gen : entity work.baudrate_gen
		port map (clk => clk, rst => rst, tick => tick);

	data <= rx_data;

	-- Registers
	process (clk, rst)
	begin
		if rst = '1' then
			state <= IDLE;
			n <= (others => '0');
			rx_data <= (others => '0');
			sample_count <= (others => '0');
		elsif rising_edge(clk) then
			state <= next_state;
			n <= next_n;
			rx_data <= next_rx_data;
			sample_count <= next_sample_count;
		end if;
	end process;

	-- Next state logic
	process (state, rx, tick, n, rx_data, sample_count)
	begin
		-- Defaults
		next_state <= state;
		next_n <= n;
		next_rx_data <= rx_data;
		next_sample_count <= sample_count;
		done <= '0';

		case state is
			when IDLE =>
				-- Start of transmission detected
				if rx = '0' then
					-- Reset sampling counter
					next_sample_count <= (others => '0');
					next_state <= START;
				end if;

			when START =>
				-- Synchronize to tick signal generated by the baudrate generator
				if tick = '1' then
					-- Wait for the middle of the start bit
					if sample_count < 7 then
						next_sample_count <= sample_count + 1;
					else
						-- Reset sampling counter, start receiving data bits
						next_sample_count <= (others => '0');
						next_state <= RDATA;
						next_n <= (others => '0');
					end if;
				end if;

			when RDATA =>
				if tick = '1' then
					-- Wait for the middle of a data bit
					if sample_count < 15 then
						next_sample_count <= sample_count + 1;
					else
						-- Reset sampling counter
						next_sample_count <= (others => '0');
						-- Sample data bit
						next_rx_data <= rx & rx_data(7 downto 1);
						-- Receive next data bit
						if n < 7 then
							next_n <= n + 1;
						else
							-- All data bits received, wait for stop bit
							next_state <= STOP;
						end if;
					end if;
				end if;

			when STOP =>
				if tick = '1' then
					-- Wait until signal becomes idle again
					if sample_count < 15 then
						next_sample_count <= sample_count + 1;
					else
						-- Jump back to idle state and indicate received data is valid
						next_state <= IDLE;
						done <= '1';
					end if;
				end if;
		end case;
	end process;
end architecture;
